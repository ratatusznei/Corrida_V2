y; ~xy  PISTA 1                       cIYTL 1 �uH�u��( ���u 